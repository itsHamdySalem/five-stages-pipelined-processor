LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY ALU IS
PORT (
X : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
Y : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
Func : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
F : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
Z : OUT STD_LOGIC; -- zero flag
N : OUT STD_LOGIC; -- negative flag
C : OUT STD_LOGIC -- carrry flag
);
END ALU;

ARCHITECTURE Behavioral OF ALU IS

BEGIN

END ARCHITECTURE;